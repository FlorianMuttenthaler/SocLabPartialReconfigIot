-------------------------------------------------------------------------------
--
-- black_white_filter_logic Testbench
--
-------------------------------------------------------------------------------
--

library ieee;
use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

use work.black_white_filter_logic_pkg.all;


--  A testbench has no ports.
entity black_white_filter_logic_tb is
end black_white_filter_logic_tb;
--
-------------------------------------------------------------------------------
--
architecture beh of black_white_filter_logic_tb is

	--  Specifies which entity is bound with the component.
	for black_white_filter_logic_0: black_white_filter_logic use entity work.black_white_filter_logic;	

	constant clk_period : time := 1 ns;
	constant DATA_WIDTH : integer := 32;
	constant THRESHOLD	: integer := 128;
	
	signal Clk : std_logic := '0';
	signal testdata1_in		:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata2_in		:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata3_in		:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata4_in		:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata1_out	:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata2_out	:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata3_out	:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata4_out	:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
begin

	--  Component instantiation.
	black_white_filter_logic_0: black_white_filter_logic
		generic map(
			C_S_AXI_DATA_WIDTH	=> DATA_WIDTH,
			THRESHOLD			=> THRESHOLD
		)
		port map (
			Clk => Clk,
			reg001in	=>	testdata1_in,
			reg002in   	=>	testdata2_in,
			reg003in   	=>	testdata3_in,
			reg004in   	=>	testdata4_in,
			reg005in   	=>	(others => '0'),
			reg006in   	=>	(others => '0'),
			reg007in   	=>	(others => '0'),
			reg008in   	=>	(others => '0'),
			reg009in   	=>	(others => '0'),
			reg010in   	=>	(others => '0'),
			reg011in   	=>	(others => '0'),
			reg012in   	=>	(others => '0'),
			reg013in   	=>	(others => '0'),
			reg014in   	=>	(others => '0'),
			reg015in   	=>	(others => '0'),
			reg016in   	=>	(others => '0'),
			reg017in   	=>	(others => '0'),
			reg018in   	=>	(others => '0'),
			reg019in   	=>	(others => '0'),
			reg020in   	=>	(others => '0'),
			reg021in   	=>	(others => '0'),
			reg022in   	=>	(others => '0'),
			reg023in   	=>	(others => '0'),
			reg024in   	=>	(others => '0'),
			reg025in   	=>	(others => '0'),
			reg026in   	=>	(others => '0'),
			reg027in   	=>	(others => '0'),
			reg028in   	=>	(others => '0'),
			reg029in   	=>	(others => '0'),
			reg030in   	=>	(others => '0'),
			reg031in   	=>	(others => '0'),
			reg032in   	=>	(others => '0'),
			reg033in   	=>	(others => '0'),
			reg034in   	=>	(others => '0'),
			reg035in   	=>	(others => '0'),
			reg036in   	=>	(others => '0'),
			reg037in   	=>	(others => '0'),
			reg038in   	=>	(others => '0'),
			reg039in   	=>	(others => '0'),
			reg040in   	=>	(others => '0'),
			reg041in   	=>	(others => '0'),
			reg042in   	=>	(others => '0'),
			reg043in   	=>	(others => '0'),
			reg044in   	=>	(others => '0'),
			reg045in   	=>	(others => '0'),
			reg046in   	=>	(others => '0'),
			reg047in   	=>	(others => '0'),
			reg048in   	=>	(others => '0'),
			reg049in   	=>	(others => '0'),
			reg050in   	=>	(others => '0'),
			reg051in   	=>	(others => '0'),
			reg052in   	=>	(others => '0'),
			reg053in   	=>	(others => '0'),
			reg054in   	=>	(others => '0'),
			reg055in   	=>	(others => '0'),
			reg056in   	=>	(others => '0'),
			reg057in   	=>	(others => '0'),
			reg058in   	=>	(others => '0'),
			reg059in   	=>	(others => '0'),
			reg060in   	=>	(others => '0'),
			reg061in   	=>	(others => '0'),
			reg062in   	=>	(others => '0'),
			reg063in   	=>	(others => '0'),
			reg064in   	=>	(others => '0'),
			reg065in   	=>	(others => '0'),
			reg066in   	=>	(others => '0'),
			reg067in   	=>	(others => '0'),
			reg068in   	=>	(others => '0'),
			reg069in   	=>	(others => '0'),
			reg070in   	=>	(others => '0'),
			reg071in   	=>	(others => '0'),
			reg072in   	=>	(others => '0'),
			reg073in   	=>	(others => '0'),
			reg074in   	=>	(others => '0'),
			reg075in   	=>	(others => '0'),
			reg076in   	=>	(others => '0'),
			reg077in   	=>	(others => '0'),
			reg078in   	=>	(others => '0'),
			reg079in   	=>	(others => '0'),
			reg080in   	=>	(others => '0'),
			reg081in   	=>	(others => '0'),
			reg082in   	=>	(others => '0'),
			reg083in   	=>	(others => '0'),
			reg084in   	=>	(others => '0'),
			reg085in   	=>	(others => '0'),
			reg086in   	=>	(others => '0'),
			reg087in   	=>	(others => '0'),
			reg088in   	=>	(others => '0'),
			reg089in   	=>	(others => '0'),
			reg090in   	=>	(others => '0'),
			reg091in   	=>	(others => '0'),
			reg092in   	=>	(others => '0'),
			reg093in   	=>	(others => '0'),
			reg094in   	=>	(others => '0'),
			reg095in   	=>	(others => '0'),
			reg096in   	=>	(others => '0'),
			reg097in   	=>	(others => '0'),
			reg098in   	=>	(others => '0'),
			reg099in   	=>	(others => '0'),
			reg100in   	=>	(others => '0'),
			reg101in   	=>	(others => '0'),
			reg102in   	=>	(others => '0'),
			reg103in   	=>	(others => '0'),
			reg104in   	=>	(others => '0'),
			reg105in   	=>	(others => '0'),
			reg106in   	=>	(others => '0'),
			reg107in   	=>	(others => '0'),
			reg108in   	=>	(others => '0'),
			reg109in   	=>	(others => '0'),
			reg110in   	=>	(others => '0'),
			reg111in   	=>	(others => '0'),
			reg112in   	=>	(others => '0'),
			reg113in   	=>	(others => '0'),
			reg114in   	=>	(others => '0'),
			reg115in   	=>	(others => '0'),
			reg116in   	=>	(others => '0'),
			reg117in   	=>	(others => '0'),
			reg118in   	=>	(others => '0'),
			reg119in   	=>	(others => '0'),
			reg120in   	=>	(others => '0'),
			reg121in   	=>	(others => '0'),
			reg122in   	=>	(others => '0'),
			reg123in   	=>	(others => '0'),
			reg124in   	=>	(others => '0'),
			reg125in   	=>	(others => '0'),
			reg126in   	=>	(others => '0'),
			reg127in   	=>	(others => '0'),
			reg128in   	=>	(others => '0'),
			reg129in   	=>	(others => '0'),
			reg130in   	=>	(others => '0'),
			reg131in   	=>	(others => '0'),
			reg132in   	=>	(others => '0'),
			reg133in   	=>	(others => '0'),
			reg134in   	=>	(others => '0'),
			reg135in   	=>	(others => '0'),
			reg136in   	=>	(others => '0'),
			reg137in   	=>	(others => '0'),
			reg138in   	=>	(others => '0'),
			reg139in   	=>	(others => '0'),
			reg140in   	=>	(others => '0'),
			reg141in   	=>	(others => '0'),
			reg142in   	=>	(others => '0'),
			reg143in   	=>	(others => '0'),
			reg144in   	=>	(others => '0'),
			reg145in   	=>	(others => '0'),
			reg146in   	=>	(others => '0'),
			reg147in   	=>	(others => '0'),
			reg148in   	=>	(others => '0'),
			reg149in   	=>	(others => '0'),
			reg150in   	=>	(others => '0'),
			reg151in   	=>	(others => '0'),
			reg152in   	=>	(others => '0'),
			reg153in   	=>	(others => '0'),
			reg154in   	=>	(others => '0'),
			reg155in   	=>	(others => '0'),
			reg156in   	=>	(others => '0'),
			reg157in   	=>	(others => '0'),
			reg158in   	=>	(others => '0'),
			reg159in   	=>	(others => '0'),
			reg160in   	=>	(others => '0'),
			reg161in   	=>	(others => '0'),
			reg162in   	=>	(others => '0'),
			reg163in   	=>	(others => '0'),
			reg164in   	=>	(others => '0'),
			reg165in   	=>	(others => '0'),
			reg166in   	=>	(others => '0'),
			reg167in   	=>	(others => '0'),
			reg168in   	=>	(others => '0'),
			reg169in   	=>	(others => '0'),
			reg170in   	=>	(others => '0'),
			reg171in   	=>	(others => '0'),
			reg172in   	=>	(others => '0'),
			reg173in   	=>	(others => '0'),
			reg174in   	=>	(others => '0'),
			reg175in   	=>	(others => '0'),
			reg176in   	=>	(others => '0'),
			reg177in   	=>	(others => '0'),
			reg178in   	=>	(others => '0'),
			reg179in   	=>	(others => '0'),
			reg180in   	=>	(others => '0'),
			reg181in   	=>	(others => '0'),
			reg182in   	=>	(others => '0'),
			reg183in   	=>	(others => '0'),
			reg184in   	=>	(others => '0'),
			reg185in   	=>	(others => '0'),
			reg186in   	=>	(others => '0'),
			reg187in   	=>	(others => '0'),
			reg188in   	=>	(others => '0'),
			reg189in   	=>	(others => '0'),
			reg190in   	=>	(others => '0'),
			reg191in   	=>	(others => '0'),
			reg192in   	=>	(others => '0'),
			reg193in   	=>	(others => '0'),
			reg194in   	=>	(others => '0'),
			reg195in   	=>	(others => '0'),
			reg196in   	=>	(others => '0'),
			reg197in   	=>	(others => '0'),
			reg198in   	=>	(others => '0'),
			reg199in   	=>	(others => '0'),
			reg200in   	=>	(others => '0'),
			reg201in   	=>	(others => '0'),
			reg202in   	=>	(others => '0'),
			reg203in   	=>	(others => '0'),
			reg204in   	=>	(others => '0'),
			reg205in   	=>	(others => '0'),
			reg206in   	=>	(others => '0'),
			reg207in   	=>	(others => '0'),
			reg208in   	=>	(others => '0'),
			reg209in   	=>	(others => '0'),
			reg210in   	=>	(others => '0'),
			reg211in   	=>	(others => '0'),
			reg212in   	=>	(others => '0'),
			reg213in   	=>	(others => '0'),
			reg214in   	=>	(others => '0'),
			reg215in   	=>	(others => '0'),
			reg216in   	=>	(others => '0'),
			reg217in   	=>	(others => '0'),
			reg218in   	=>	(others => '0'),
			reg219in   	=>	(others => '0'),
			reg220in   	=>	(others => '0'),
			reg221in   	=>	(others => '0'),
			reg222in   	=>	(others => '0'),
			reg223in   	=>	(others => '0'),
			reg224in   	=>	(others => '0'),
			reg225in   	=>	(others => '0'),
			reg226in   	=>	(others => '0'),
			reg227in   	=>	(others => '0'),
			reg228in   	=>	(others => '0'),
			reg229in   	=>	(others => '0'),
			reg230in   	=>	(others => '0'),
			reg231in   	=>	(others => '0'),
			reg232in   	=>	(others => '0'),
			reg233in   	=>	(others => '0'),
			reg234in   	=>	(others => '0'),
			reg235in   	=>	(others => '0'),
			reg236in   	=>	(others => '0'),
			reg237in   	=>	(others => '0'),
			reg238in   	=>	(others => '0'),
			reg239in   	=>	(others => '0'),
			reg240in   	=>	(others => '0'),
			reg241in   	=>	(others => '0'),
			reg242in   	=>	(others => '0'),
			reg243in   	=>	(others => '0'),
			reg244in   	=>	(others => '0'),
			reg245in   	=>	(others => '0'),
			reg246in   	=>	(others => '0'),
			reg247in   	=>	(others => '0'),
			reg248in   	=>	(others => '0'),
			reg249in   	=>	(others => '0'),
			reg250in   	=>	(others => '0'),
			reg251in   	=>	(others => '0'),
			reg252in   	=>	(others => '0'),
			reg253in   	=>	(others => '0'),
			reg254in   	=>	(others => '0'),
			reg255in   	=>	(others => '0'),
			reg256in   	=>	(others => '0'),
			reg001out   =>	testdata1_out,
			reg002out   =>	testdata2_out,
			reg003out   =>	testdata3_out,
			reg004out   =>	testdata4_out,
			reg005out   =>	(others => '0'),
			reg006out   =>	(others => '0'),
			reg007out   =>	(others => '0'),
			reg008out   =>	(others => '0'),
			reg009out   =>	(others => '0'),
			reg010out   =>	(others => '0'),
			reg011out   =>	(others => '0'),
			reg012out   =>	(others => '0'),
			reg013out   =>	(others => '0'),
			reg014out   =>	(others => '0'),
			reg015out   =>	(others => '0'),
			reg016out   =>	(others => '0'),
			reg017out   =>	(others => '0'),
			reg018out   =>	(others => '0'),
			reg019out   =>	(others => '0'),
			reg020out   =>	(others => '0'),
			reg021out   =>	(others => '0'),
			reg022out   =>	(others => '0'),
			reg023out   =>	(others => '0'),
			reg024out   =>	(others => '0'),
			reg025out   =>	(others => '0'),
			reg026out   =>	(others => '0'),
			reg027out   =>	(others => '0'),
			reg028out   =>	(others => '0'),
			reg029out   =>	(others => '0'),
			reg030out   =>	(others => '0'),
			reg031out   =>	(others => '0'),
			reg032out   =>	(others => '0'),
			reg033out   =>	(others => '0'),
			reg034out   =>	(others => '0'),
			reg035out   =>	(others => '0'),
			reg036out   =>	(others => '0'),
			reg037out   =>	(others => '0'),
			reg038out   =>	(others => '0'),
			reg039out   =>	(others => '0'),
			reg040out   =>	(others => '0'),
			reg041out   =>	(others => '0'),
			reg042out   =>	(others => '0'),
			reg043out   =>	(others => '0'),
			reg044out   =>	(others => '0'),
			reg045out   =>	(others => '0'),
			reg046out   =>	(others => '0'),
			reg047out   =>	(others => '0'),
			reg048out   =>	(others => '0'),
			reg049out   =>	(others => '0'),
			reg050out   =>	(others => '0'),
			reg051out   =>	(others => '0'),
			reg052out   =>	(others => '0'),
			reg053out   =>	(others => '0'),
			reg054out   =>	(others => '0'),
			reg055out   =>	(others => '0'),
			reg056out   =>	(others => '0'),
			reg057out   =>	(others => '0'),
			reg058out   =>	(others => '0'),
			reg059out   =>	(others => '0'),
			reg060out   =>	(others => '0'),
			reg061out   =>	(others => '0'),
			reg062out   =>	(others => '0'),
			reg063out   =>	(others => '0'),
			reg064out   =>	(others => '0'),
			reg065out   =>	(others => '0'),
			reg066out   =>	(others => '0'),
			reg067out   =>	(others => '0'),
			reg068out   =>	(others => '0'),
			reg069out   =>	(others => '0'),
			reg070out   =>	(others => '0'),
			reg071out   =>	(others => '0'),
			reg072out   =>	(others => '0'),
			reg073out   =>	(others => '0'),
			reg074out   =>	(others => '0'),
			reg075out   =>	(others => '0'),
			reg076out   =>	(others => '0'),
			reg077out   =>	(others => '0'),
			reg078out   =>	(others => '0'),
			reg079out   =>	(others => '0'),
			reg080out   =>	(others => '0'),
			reg081out   =>	(others => '0'),
			reg082out   =>	(others => '0'),
			reg083out   =>	(others => '0'),
			reg084out   =>	(others => '0'),
			reg085out   =>	(others => '0'),
			reg086out   =>	(others => '0'),
			reg087out   =>	(others => '0'),
			reg088out   =>	(others => '0'),
			reg089out   =>	(others => '0'),
			reg090out   =>	(others => '0'),
			reg091out   =>	(others => '0'),
			reg092out   =>	(others => '0'),
			reg093out   =>	(others => '0'),
			reg094out   =>	(others => '0'),
			reg095out   =>	(others => '0'),
			reg096out   =>	(others => '0'),
			reg097out   =>	(others => '0'),
			reg098out   =>	(others => '0'),
			reg099out   =>	(others => '0'),
			reg100out   =>	(others => '0'),
			reg101out   =>	(others => '0'),
			reg102out   =>	(others => '0'),
			reg103out   =>	(others => '0'),
			reg104out   =>	(others => '0'),
			reg105out   =>	(others => '0'),
			reg106out   =>	(others => '0'),
			reg107out   =>	(others => '0'),
			reg108out   =>	(others => '0'),
			reg109out   =>	(others => '0'),
			reg110out   =>	(others => '0'),
			reg111out   =>	(others => '0'),
			reg112out   =>	(others => '0'),
			reg113out   =>	(others => '0'),
			reg114out   =>	(others => '0'),
			reg115out   =>	(others => '0'),
			reg116out   =>	(others => '0'),
			reg117out   =>	(others => '0'),
			reg118out   =>	(others => '0'),
			reg119out   =>	(others => '0'),
			reg120out   =>	(others => '0'),
			reg121out   =>	(others => '0'),
			reg122out   =>	(others => '0'),
			reg123out   =>	(others => '0'),
			reg124out   =>	(others => '0'),
			reg125out   =>	(others => '0'),
			reg126out   =>	(others => '0'),
			reg127out   =>	(others => '0'),
			reg128out   =>	(others => '0'),
			reg129out   =>	(others => '0'),
			reg130out   =>	(others => '0'),
			reg131out   =>	(others => '0'),
			reg132out   =>	(others => '0'),
			reg133out   =>	(others => '0'),
			reg134out   =>	(others => '0'),
			reg135out   =>	(others => '0'),
			reg136out   =>	(others => '0'),
			reg137out   =>	(others => '0'),
			reg138out   =>	(others => '0'),
			reg139out   =>	(others => '0'),
			reg140out   =>	(others => '0'),
			reg141out   =>	(others => '0'),
			reg142out   =>	(others => '0'),
			reg143out   =>	(others => '0'),
			reg144out   =>	(others => '0'),
			reg145out   =>	(others => '0'),
			reg146out   =>	(others => '0'),
			reg147out   =>	(others => '0'),
			reg148out   =>	(others => '0'),
			reg149out   =>	(others => '0'),
			reg150out   =>	(others => '0'),
			reg151out   =>	(others => '0'),
			reg152out   =>	(others => '0'),
			reg153out   =>	(others => '0'),
			reg154out   =>	(others => '0'),
			reg155out   =>	(others => '0'),
			reg156out   =>	(others => '0'),
			reg157out   =>	(others => '0'),
			reg158out   =>	(others => '0'),
			reg159out   =>	(others => '0'),
			reg160out   =>	(others => '0'),
			reg161out   =>	(others => '0'),
			reg162out   =>	(others => '0'),
			reg163out   =>	(others => '0'),
			reg164out   =>	(others => '0'),
			reg165out   =>	(others => '0'),
			reg166out   =>	(others => '0'),
			reg167out   =>	(others => '0'),
			reg168out   =>	(others => '0'),
			reg169out   =>	(others => '0'),
			reg170out   =>	(others => '0'),
			reg171out   =>	(others => '0'),
			reg172out   =>	(others => '0'),
			reg173out   =>	(others => '0'),
			reg174out   =>	(others => '0'),
			reg175out   =>	(others => '0'),
			reg176out   =>	(others => '0'),
			reg177out   =>	(others => '0'),
			reg178out   =>	(others => '0'),
			reg179out   =>	(others => '0'),
			reg180out   =>	(others => '0'),
			reg181out   =>	(others => '0'),
			reg182out   =>	(others => '0'),
			reg183out   =>	(others => '0'),
			reg184out   =>	(others => '0'),
			reg185out   =>	(others => '0'),
			reg186out   =>	(others => '0'),
			reg187out   =>	(others => '0'),
			reg188out   =>	(others => '0'),
			reg189out   =>	(others => '0'),
			reg190out   =>	(others => '0'),
			reg191out   =>	(others => '0'),
			reg192out   =>	(others => '0'),
			reg193out   =>	(others => '0'),
			reg194out   =>	(others => '0'),
			reg195out   =>	(others => '0'),
			reg196out   =>	(others => '0'),
			reg197out   =>	(others => '0'),
			reg198out   =>	(others => '0'),
			reg199out   =>	(others => '0'),
			reg200out   =>	(others => '0'),
			reg201out   =>	(others => '0'),
			reg202out   =>	(others => '0'),
			reg203out   =>	(others => '0'),
			reg204out   =>	(others => '0'),
			reg205out   =>	(others => '0'),
			reg206out   =>	(others => '0'),
			reg207out   =>	(others => '0'),
			reg208out   =>	(others => '0'),
			reg209out   =>	(others => '0'),
			reg210out   =>	(others => '0'),
			reg211out   =>	(others => '0'),
			reg212out   =>	(others => '0'),
			reg213out   =>	(others => '0'),
			reg214out   =>	(others => '0'),
			reg215out   =>	(others => '0'),
			reg216out   =>	(others => '0'),
			reg217out   =>	(others => '0'),
			reg218out   =>	(others => '0'),
			reg219out   =>	(others => '0'),
			reg220out   =>	(others => '0'),
			reg221out   =>	(others => '0'),
			reg222out   =>	(others => '0'),
			reg223out   =>	(others => '0'),
			reg224out   =>	(others => '0'),
			reg225out   =>	(others => '0'),
			reg226out   =>	(others => '0'),
			reg227out   =>	(others => '0'),
			reg228out   =>	(others => '0'),
			reg229out   =>	(others => '0'),
			reg230out   =>	(others => '0'),
			reg231out   =>	(others => '0'),
			reg232out   =>	(others => '0'),
			reg233out   =>	(others => '0'),
			reg234out   =>	(others => '0'),
			reg235out   =>	(others => '0'),
			reg236out   =>	(others => '0'),
			reg237out   =>	(others => '0'),
			reg238out   =>	(others => '0'),
			reg239out   =>	(others => '0'),
			reg240out   =>	(others => '0'),
			reg241out   =>	(others => '0'),
			reg242out   =>	(others => '0'),
			reg243out   =>	(others => '0'),
			reg244out   =>	(others => '0'),
			reg245out   =>	(others => '0'),
			reg246out   =>	(others => '0'),
			reg247out   =>	(others => '0'),
			reg248out   =>	(others => '0'),
			reg249out   =>	(others => '0'),
			reg250out   =>	(others => '0'),
			reg251out   =>	(others => '0'),
			reg252out   =>	(others => '0'),
			reg253out   =>	(others => '0'),
			reg254out   =>	(others => '0'),
			reg255out   =>	(others => '0'),
			reg256out   =>	(others => '0')
		);
		
	Clk_process : process
	
	begin
		Clk <= '0';
		wait for clk_period/2;
		Clk <= '1';
		wait for clk_period/2;

	end process clk_process;	

	--  This process does the real job.
	stimuli : process

	begin

		wait for 10 ns;

		testdata2_in <= (others => '1');
		
		wait for 2 ns;
		
		--assert testdata2_out = "11111111111111111111111111111111" report "Test data 2 correct" severity note;
		
		wait for 2 ns;
			
		testdata3_in <= "00000000000000000000000010000000";
		
		wait for 2 ns;
		
		--assert testdata3_out = "11111111111111111111111111111111" report "Test data 3 correct" severity note;
		
		wait for 2 ns;

		testdata4_in <= "00000000000000000000000001111111";
		
		wait for 2 ns;
		
		--assert testdata4_out = "00000000000000000000000000000000" report "Test data 4 correct" severity note;
		
		wait for 2 ns;
		
		testdata1_in <= (others => '0');
		
		wait for 2 ns;
		
		--assert testdata1_out = "00000000000000000000000000000000" report "Test data 1 correct" severity note;
		
		wait for 2 ns;
		
		assert false report "end of test" severity note;

		--  Wait forever; this will finish the simulation.
		wait;

	end process stimuli;

end beh;
--
-------------------------------------------------------------------------------
