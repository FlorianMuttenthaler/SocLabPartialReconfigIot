-------------------------------------------------------------------------------
--
-- black_white_filter_logic Testbench
--
-------------------------------------------------------------------------------
--

library ieee;
use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

use work.black_white_filter_logic_pkg.all;


--  A testbench has no ports.
entity black_white_filter_logic_tb is
end black_white_filter_logic_tb;
--
-------------------------------------------------------------------------------
--
architecture beh of black_white_filter_logic_tb is

	--  Specifies which entity is bound with the component.
	for black_white_filter_logic_0: black_white_filter_logic use entity work.black_white_filter_logic;	

	constant clk_period : time := 1 ns;
	constant DATA_WIDTH : integer := 32;
	constant THRESHOLD	: integer := 128;
	
	signal Clk : std_logic := '0';
	signal testdata1_in		:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata2_in		:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata3_in		:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata4_in		:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata1_out	:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata2_out	:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata3_out	:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
	signal testdata4_out	:	std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
begin

	--  Component instantiation.
	black_white_filter_logic_0: black_white_filter_logic
		generic map(
			C_S_AXI_DATA_WIDTH	=> DATA_WIDTH,
			THRESHOLD			=> THRESHOLD
		)
		port map (
			Clk => Clk,
			reg001in	=>	testdata1_in,
			reg002in   	=>	testdata2_in,
			reg003in   	=>	testdata3_in,
			reg004in   	=>	testdata4_in,
			reg005in   	=>	(others => '0'),
			reg006in   	=>	(others => '0'),
			reg007in   	=>	(others => '0'),
			reg008in   	=>	(others => '0'),
			reg009in   	=>	(others => '0'),
			reg010in   	=>	(others => '0'),
			reg011in   	=>	(others => '0'),
			reg012in   	=>	(others => '0'),
			reg013in   	=>	(others => '0'),
			reg014in   	=>	(others => '0'),
			reg015in   	=>	(others => '0'),
			reg016in   	=>	(others => '0'),
			reg017in   	=>	(others => '0'),
			reg018in   	=>	(others => '0'),
			reg019in   	=>	(others => '0'),
			reg020in   	=>	(others => '0'),
			reg021in   	=>	(others => '0'),
			reg022in   	=>	(others => '0'),
			reg023in   	=>	(others => '0'),
			reg024in   	=>	(others => '0'),
			reg025in   	=>	(others => '0'),
			reg026in   	=>	(others => '0'),
			reg027in   	=>	(others => '0'),
			reg028in   	=>	(others => '0'),
			reg029in   	=>	(others => '0'),
			reg030in   	=>	(others => '0'),
			reg031in   	=>	(others => '0'),
			reg032in   	=>	(others => '0'),
			reg033in   	=>	(others => '0'),
			reg034in   	=>	(others => '0'),
			reg035in   	=>	(others => '0'),
			reg036in   	=>	(others => '0'),
			reg037in   	=>	(others => '0'),
			reg038in   	=>	(others => '0'),
			reg039in   	=>	(others => '0'),
			reg040in   	=>	(others => '0'),
			reg041in   	=>	(others => '0'),
			reg042in   	=>	(others => '0'),
			reg043in   	=>	(others => '0'),
			reg044in   	=>	(others => '0'),
			reg045in   	=>	(others => '0'),
			reg046in   	=>	(others => '0'),
			reg047in   	=>	(others => '0'),
			reg048in   	=>	(others => '0'),
			reg049in   	=>	(others => '0'),
			reg050in   	=>	(others => '0'),
			reg051in   	=>	(others => '0'),
			reg052in   	=>	(others => '0'),
			reg053in   	=>	(others => '0'),
			reg054in   	=>	(others => '0'),
			reg055in   	=>	(others => '0'),
			reg056in   	=>	(others => '0'),
			reg057in   	=>	(others => '0'),
			reg058in   	=>	(others => '0'),
			reg059in   	=>	(others => '0'),
			reg060in   	=>	(others => '0'),
			reg061in   	=>	(others => '0'),
			reg062in   	=>	(others => '0'),
			reg063in   	=>	(others => '0'),
			reg064in   	=>	(others => '0'),
			reg065in   	=>	(others => '0'),
			reg066in   	=>	(others => '0'),
			reg067in   	=>	(others => '0'),
			reg068in   	=>	(others => '0'),
			reg069in   	=>	(others => '0'),
			reg070in   	=>	(others => '0'),
			reg071in   	=>	(others => '0'),
			reg072in   	=>	(others => '0'),
			reg073in   	=>	(others => '0'),
			reg074in   	=>	(others => '0'),
			reg075in   	=>	(others => '0'),
			reg076in   	=>	(others => '0'),
			reg077in   	=>	(others => '0'),
			reg078in   	=>	(others => '0'),
			reg079in   	=>	(others => '0'),
			reg080in   	=>	(others => '0'),
			reg081in   	=>	(others => '0'),
			reg082in   	=>	(others => '0'),
			reg083in   	=>	(others => '0'),
			reg084in   	=>	(others => '0'),
			reg085in   	=>	(others => '0'),
			reg086in   	=>	(others => '0'),
			reg087in   	=>	(others => '0'),
			reg088in   	=>	(others => '0'),
			reg089in   	=>	(others => '0'),
			reg090in   	=>	(others => '0'),
			reg091in   	=>	(others => '0'),
			reg092in   	=>	(others => '0'),
			reg093in   	=>	(others => '0'),
			reg094in   	=>	(others => '0'),
			reg095in   	=>	(others => '0'),
			reg096in   	=>	(others => '0'),
			reg097in   	=>	(others => '0'),
			reg098in   	=>	(others => '0'),
			reg099in   	=>	(others => '0'),
			reg100in   	=>	(others => '0'),
			reg101in   	=>	(others => '0'),
			reg102in   	=>	(others => '0'),
			reg103in   	=>	(others => '0'),
			reg104in   	=>	(others => '0'),
			reg105in   	=>	(others => '0'),
			reg106in   	=>	(others => '0'),
			reg107in   	=>	(others => '0'),
			reg108in   	=>	(others => '0'),
			reg109in   	=>	(others => '0'),
			reg110in   	=>	(others => '0'),
			reg111in   	=>	(others => '0'),
			reg112in   	=>	(others => '0'),
			reg113in   	=>	(others => '0'),
			reg114in   	=>	(others => '0'),
			reg115in   	=>	(others => '0'),
			reg116in   	=>	(others => '0'),
			reg117in   	=>	(others => '0'),
			reg118in   	=>	(others => '0'),
			reg119in   	=>	(others => '0'),
			reg120in   	=>	(others => '0'),
			reg121in   	=>	(others => '0'),
			reg122in   	=>	(others => '0'),
			reg123in   	=>	(others => '0'),
			reg124in   	=>	(others => '0'),
			reg125in   	=>	(others => '0'),
			reg126in   	=>	(others => '0'),
			reg127in   	=>	(others => '0'),
			reg128in   	=>	(others => '0'),
			reg129in   	=>	(others => '0'),
			reg130in   	=>	(others => '0'),
			reg131in   	=>	(others => '0'),
			reg132in   	=>	(others => '0'),
			reg133in   	=>	(others => '0'),
			reg134in   	=>	(others => '0'),
			reg135in   	=>	(others => '0'),
			reg136in   	=>	(others => '0'),
			reg137in   	=>	(others => '0'),
			reg138in   	=>	(others => '0'),
			reg139in   	=>	(others => '0'),
			reg140in   	=>	(others => '0'),
			reg141in   	=>	(others => '0'),
			reg142in   	=>	(others => '0'),
			reg143in   	=>	(others => '0'),
			reg144in   	=>	(others => '0'),
			reg145in   	=>	(others => '0'),
			reg146in   	=>	(others => '0'),
			reg147in   	=>	(others => '0'),
			reg148in   	=>	(others => '0'),
			reg149in   	=>	(others => '0'),
			reg150in   	=>	(others => '0'),
			reg151in   	=>	(others => '0'),
			reg152in   	=>	(others => '0'),
			reg153in   	=>	(others => '0'),
			reg154in   	=>	(others => '0'),
			reg155in   	=>	(others => '0'),
			reg156in   	=>	(others => '0'),
			reg157in   	=>	(others => '0'),
			reg158in   	=>	(others => '0'),
			reg159in   	=>	(others => '0'),
			reg160in   	=>	(others => '0'),
			reg161in   	=>	(others => '0'),
			reg162in   	=>	(others => '0'),
			reg163in   	=>	(others => '0'),
			reg164in   	=>	(others => '0'),
			reg165in   	=>	(others => '0'),
			reg166in   	=>	(others => '0'),
			reg167in   	=>	(others => '0'),
			reg168in   	=>	(others => '0'),
			reg169in   	=>	(others => '0'),
			reg170in   	=>	(others => '0'),
			reg171in   	=>	(others => '0'),
			reg172in   	=>	(others => '0'),
			reg173in   	=>	(others => '0'),
			reg174in   	=>	(others => '0'),
			reg175in   	=>	(others => '0'),
			reg176in   	=>	(others => '0'),
			reg177in   	=>	(others => '0'),
			reg178in   	=>	(others => '0'),
			reg179in   	=>	(others => '0'),
			reg180in   	=>	(others => '0'),
			reg181in   	=>	(others => '0'),
			reg182in   	=>	(others => '0'),
			reg183in   	=>	(others => '0'),
			reg184in   	=>	(others => '0'),
			reg185in   	=>	(others => '0'),
			reg186in   	=>	(others => '0'),
			reg187in   	=>	(others => '0'),
			reg188in   	=>	(others => '0'),
			reg189in   	=>	(others => '0'),
			reg190in   	=>	(others => '0'),
			reg191in   	=>	(others => '0'),
			reg192in   	=>	(others => '0'),
			reg193in   	=>	(others => '0'),
			reg194in   	=>	(others => '0'),
			reg195in   	=>	(others => '0'),
			reg196in   	=>	(others => '0'),
			reg197in   	=>	(others => '0'),
			reg198in   	=>	(others => '0'),
			reg199in   	=>	(others => '0'),
			reg200in   	=>	(others => '0'),
			reg201in   	=>	(others => '0'),
			reg202in   	=>	(others => '0'),
			reg203in   	=>	(others => '0'),
			reg204in   	=>	(others => '0'),
			reg205in   	=>	(others => '0'),
			reg206in   	=>	(others => '0'),
			reg207in   	=>	(others => '0'),
			reg208in   	=>	(others => '0'),
			reg209in   	=>	(others => '0'),
			reg210in   	=>	(others => '0'),
			reg211in   	=>	(others => '0'),
			reg212in   	=>	(others => '0'),
			reg213in   	=>	(others => '0'),
			reg214in   	=>	(others => '0'),
			reg215in   	=>	(others => '0'),
			reg216in   	=>	(others => '0'),
			reg217in   	=>	(others => '0'),
			reg218in   	=>	(others => '0'),
			reg219in   	=>	(others => '0'),
			reg220in   	=>	(others => '0'),
			reg221in   	=>	(others => '0'),
			reg222in   	=>	(others => '0'),
			reg223in   	=>	(others => '0'),
			reg224in   	=>	(others => '0'),
			reg225in   	=>	(others => '0'),
			reg226in   	=>	(others => '0'),
			reg227in   	=>	(others => '0'),
			reg228in   	=>	(others => '0'),
			reg229in   	=>	(others => '0'),
			reg230in   	=>	(others => '0'),
			reg231in   	=>	(others => '0'),
			reg232in   	=>	(others => '0'),
			reg233in   	=>	(others => '0'),
			reg234in   	=>	(others => '0'),
			reg235in   	=>	(others => '0'),
			reg236in   	=>	(others => '0'),
			reg237in   	=>	(others => '0'),
			reg238in   	=>	(others => '0'),
			reg239in   	=>	(others => '0'),
			reg240in   	=>	(others => '0'),
			reg241in   	=>	(others => '0'),
			reg242in   	=>	(others => '0'),
			reg243in   	=>	(others => '0'),
			reg244in   	=>	(others => '0'),
			reg245in   	=>	(others => '0'),
			reg246in   	=>	(others => '0'),
			reg247in   	=>	(others => '0'),
			reg248in   	=>	(others => '0'),
			reg249in   	=>	(others => '0'),
			reg250in   	=>	(others => '0'),
			reg251in   	=>	(others => '0'),
			reg252in   	=>	(others => '0'),
			reg253in   	=>	(others => '0'),
			reg254in   	=>	(others => '0'),
			reg255in   	=>	(others => '0'),
			reg256in   	=>	(others => '0'),
			reg001out   =>	testdata1_out,
			reg002out   =>	testdata2_out,
			reg003out   =>	testdata3_out,
			reg004out   =>	testdata4_out,
			reg005out   =>	open,
			reg006out   =>	open,
			reg007out   =>	open,
			reg008out   =>	open,
			reg009out   =>	open,
			reg010out   =>	open,
			reg011out   =>	open,
			reg012out   =>	open,
			reg013out   =>	open,
			reg014out   =>	open,
			reg015out   =>	open,
			reg016out   =>	open,
			reg017out   =>	open,
			reg018out   =>	open,
			reg019out   =>	open,
			reg020out   =>	open,
			reg021out   =>	open,
			reg022out   =>	open,
			reg023out   =>	open,
			reg024out   =>	open,
			reg025out   =>	open,
			reg026out   =>	open,
			reg027out   =>	open,
			reg028out   =>	open,
			reg029out   =>	open,
			reg030out   =>	open,
			reg031out   =>	open,
			reg032out   =>	open,
			reg033out   =>	open,
			reg034out   =>	open,
			reg035out   =>	open,
			reg036out   =>	open,
			reg037out   =>	open,
			reg038out   =>	open,
			reg039out   =>	open,
			reg040out   =>	open,
			reg041out   =>	open,
			reg042out   =>	open,
			reg043out   =>	open,
			reg044out   =>	open,
			reg045out   =>	open,
			reg046out   =>	open,
			reg047out   =>	open,
			reg048out   =>	open,
			reg049out   =>	open,
			reg050out   =>	open,
			reg051out   =>	open,
			reg052out   =>	open,
			reg053out   =>	open,
			reg054out   =>	open,
			reg055out   =>	open,
			reg056out   =>	open,
			reg057out   =>	open,
			reg058out   =>	open,
			reg059out   =>	open,
			reg060out   =>	open,
			reg061out   =>	open,
			reg062out   =>	open,
			reg063out   =>	open,
			reg064out   =>	open,
			reg065out   =>	open,
			reg066out   =>	open,
			reg067out   =>	open,
			reg068out   =>	open,
			reg069out   =>	open,
			reg070out   =>	open,
			reg071out   =>	open,
			reg072out   =>	open,
			reg073out   =>	open,
			reg074out   =>	open,
			reg075out   =>	open,
			reg076out   =>	open,
			reg077out   =>	open,
			reg078out   =>	open,
			reg079out   =>	open,
			reg080out   =>	open,
			reg081out   =>	open,
			reg082out   =>	open,
			reg083out   =>	open,
			reg084out   =>	open,
			reg085out   =>	open,
			reg086out   =>	open,
			reg087out   =>	open,
			reg088out   =>	open,
			reg089out   =>	open,
			reg090out   =>	open,
			reg091out   =>	open,
			reg092out   =>	open,
			reg093out   =>	open,
			reg094out   =>	open,
			reg095out   =>	open,
			reg096out   =>	open,
			reg097out   =>	open,
			reg098out   =>	open,
			reg099out   =>	open,
			reg100out   =>	open,
			reg101out   =>	open,
			reg102out   =>	open,
			reg103out   =>	open,
			reg104out   =>	open,
			reg105out   =>	open,
			reg106out   =>	open,
			reg107out   =>	open,
			reg108out   =>	open,
			reg109out   =>	open,
			reg110out   =>	open,
			reg111out   =>	open,
			reg112out   =>	open,
			reg113out   =>	open,
			reg114out   =>	open,
			reg115out   =>	open,
			reg116out   =>	open,
			reg117out   =>	open,
			reg118out   =>	open,
			reg119out   =>	open,
			reg120out   =>	open,
			reg121out   =>	open,
			reg122out   =>	open,
			reg123out   =>	open,
			reg124out   =>	open,
			reg125out   =>	open,
			reg126out   =>	open,
			reg127out   =>	open,
			reg128out   =>	open,
			reg129out   =>	open,
			reg130out   =>	open,
			reg131out   =>	open,
			reg132out   =>	open,
			reg133out   =>	open,
			reg134out   =>	open,
			reg135out   =>	open,
			reg136out   =>	open,
			reg137out   =>	open,
			reg138out   =>	open,
			reg139out   =>	open,
			reg140out   =>	open,
			reg141out   =>	open,
			reg142out   =>	open,
			reg143out   =>	open,
			reg144out   =>	open,
			reg145out   =>	open,
			reg146out   =>	open,
			reg147out   =>	open,
			reg148out   =>	open,
			reg149out   =>	open,
			reg150out   =>	open,
			reg151out   =>	open,
			reg152out   =>	open,
			reg153out   =>	open,
			reg154out   =>	open,
			reg155out   =>	open,
			reg156out   =>	open,
			reg157out   =>	open,
			reg158out   =>	open,
			reg159out   =>	open,
			reg160out   =>	open,
			reg161out   =>	open,
			reg162out   =>	open,
			reg163out   =>	open,
			reg164out   =>	open,
			reg165out   =>	open,
			reg166out   =>	open,
			reg167out   =>	open,
			reg168out   =>	open,
			reg169out   =>	open,
			reg170out   =>	open,
			reg171out   =>	open,
			reg172out   =>	open,
			reg173out   =>	open,
			reg174out   =>	open,
			reg175out   =>	open,
			reg176out   =>	open,
			reg177out   =>	open,
			reg178out   =>	open,
			reg179out   =>	open,
			reg180out   =>	open,
			reg181out   =>	open,
			reg182out   =>	open,
			reg183out   =>	open,
			reg184out   =>	open,
			reg185out   =>	open,
			reg186out   =>	open,
			reg187out   =>	open,
			reg188out   =>	open,
			reg189out   =>	open,
			reg190out   =>	open,
			reg191out   =>	open,
			reg192out   =>	open,
			reg193out   =>	open,
			reg194out   =>	open,
			reg195out   =>	open,
			reg196out   =>	open,
			reg197out   =>	open,
			reg198out   =>	open,
			reg199out   =>	open,
			reg200out   =>	open,
			reg201out   =>	open,
			reg202out   =>	open,
			reg203out   =>	open,
			reg204out   =>	open,
			reg205out   =>	open,
			reg206out   =>	open,
			reg207out   =>	open,
			reg208out   =>	open,
			reg209out   =>	open,
			reg210out   =>	open,
			reg211out   =>	open,
			reg212out   =>	open,
			reg213out   =>	open,
			reg214out   =>	open,
			reg215out   =>	open,
			reg216out   =>	open,
			reg217out   =>	open,
			reg218out   =>	open,
			reg219out   =>	open,
			reg220out   =>	open,
			reg221out   =>	open,
			reg222out   =>	open,
			reg223out   =>	open,
			reg224out   =>	open,
			reg225out   =>	open,
			reg226out   =>	open,
			reg227out   =>	open,
			reg228out   =>	open,
			reg229out   =>	open,
			reg230out   =>	open,
			reg231out   =>	open,
			reg232out   =>	open,
			reg233out   =>	open,
			reg234out   =>	open,
			reg235out   =>	open,
			reg236out   =>	open,
			reg237out   =>	open,
			reg238out   =>	open,
			reg239out   =>	open,
			reg240out   =>	open,
			reg241out   =>	open,
			reg242out   =>	open,
			reg243out   =>	open,
			reg244out   =>	open,
			reg245out   =>	open,
			reg246out   =>	open,
			reg247out   =>	open,
			reg248out   =>	open,
			reg249out   =>	open,
			reg250out   =>	open,
			reg251out   =>	open,
			reg252out   =>	open,
			reg253out   =>	open,
			reg254out   =>	open,
			reg255out   =>	open,
			reg256out   =>	open
		);
		
	Clk_process : process
	
	begin
		Clk <= '0';
		wait for clk_period/2;
		Clk <= '1';
		wait for clk_period/2;

	end process clk_process;	

	--  This process does the real job.
	stimuli : process

	begin

		wait for 10 ns;

		testdata2_in <= (others => '1');
		
		wait for 2 ns;
		
		--assert testdata2_out = "11111111111111111111111111111111" report "Test data 2 correct" severity note;
		
		wait for 2 ns;
			
		testdata3_in <= "00000000000000000000000010000000";
		
		wait for 2 ns;
		
		--assert testdata3_out = "11111111111111111111111111111111" report "Test data 3 correct" severity note;
		
		wait for 2 ns;

		testdata4_in <= "00000000000000000000000001111111";
		
		wait for 2 ns;
		
		--assert testdata4_out = "00000000000000000000000000000000" report "Test data 4 correct" severity note;
		
		wait for 2 ns;
		
		testdata1_in <= (others => '0');
		
		wait for 2 ns;
		
		--assert testdata1_out = "00000000000000000000000000000000" report "Test data 1 correct" severity note;
		
		wait for 2 ns;
		
		assert false report "end of test" severity note;

		--  Wait forever; this will finish the simulation.
		wait;

	end process stimuli;

end beh;
--
-------------------------------------------------------------------------------
