library ieee;
use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity black_white_filter_logic is
  generic(
    -- Width of S_AXI data bus
    C_S_AXI_DATA_WIDTH	: integer	:= 32;
	THRESHOLD			: integer	:= 128
  );
  port(
    clk 	: in std_logic;
    reg001in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg002in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg003in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg004in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg005in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg006in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg007in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg008in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg009in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg010in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg011in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg012in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg013in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg014in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg015in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg016in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg017in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg018in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg019in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg020in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg021in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg022in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg023in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg024in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg025in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg026in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg027in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg028in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg029in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg030in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg031in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg032in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg033in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg034in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg035in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg036in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg037in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg038in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg039in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg040in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg041in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg042in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg043in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg044in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg045in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg046in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg047in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg048in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg049in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg050in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg051in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg052in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg053in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg054in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg055in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg056in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg057in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg058in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg059in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg060in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg061in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg062in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg063in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg064in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg065in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg066in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg067in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg068in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg069in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg070in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg071in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg072in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg073in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg074in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg075in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg076in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg077in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg078in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg079in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg080in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg081in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg082in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg083in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg084in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg085in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg086in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg087in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg088in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg089in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg090in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg091in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg092in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg093in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg094in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg095in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg096in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg097in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg098in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg099in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg100in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg101in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg102in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg103in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg104in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg105in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg106in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg107in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg108in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg109in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg110in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg111in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg112in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg113in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg114in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg115in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg116in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg117in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg118in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg119in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg120in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg121in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg122in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg123in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg124in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg125in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg126in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg127in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg128in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg129in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg130in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg131in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg132in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg133in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg134in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg135in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg136in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg137in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg138in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg139in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg140in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg141in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg142in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg143in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg144in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg145in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg146in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg147in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg148in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg149in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg150in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg151in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg152in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg153in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg154in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg155in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg156in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg157in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg158in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg159in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg160in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg161in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg162in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg163in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg164in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg165in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg166in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg167in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg168in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg169in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg170in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg171in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg172in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg173in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg174in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg175in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg176in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg177in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg178in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg179in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg180in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg181in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg182in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg183in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg184in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg185in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg186in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg187in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg188in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg189in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg190in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg191in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg192in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg193in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg194in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg195in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg196in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg197in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg198in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg199in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg200in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg201in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg202in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg203in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg204in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg205in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg206in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg207in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg208in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg209in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg210in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg211in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg212in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg213in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg214in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg215in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg216in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg217in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg218in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg219in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg220in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg221in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg222in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg223in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg224in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg225in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg226in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg227in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg228in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg229in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg230in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg231in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg232in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg233in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg234in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg235in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg236in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg237in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg238in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg239in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg240in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg241in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg242in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg243in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg244in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg245in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg246in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg247in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg248in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg249in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg250in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg251in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg252in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg253in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg254in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg255in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg256in   	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg001out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg002out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg003out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg004out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg005out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg006out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg007out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg008out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg009out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg010out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg011out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg012out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg013out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg014out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg015out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg016out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg017out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg018out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg019out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg020out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg021out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg022out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg023out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg024out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg025out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg026out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg027out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg028out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg029out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg030out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg031out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg032out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg033out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg034out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg035out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg036out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg037out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg038out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg039out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg040out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg041out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg042out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg043out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg044out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg045out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg046out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg047out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg048out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg049out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg050out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg051out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg052out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg053out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg054out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg055out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg056out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg057out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg058out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg059out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg060out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg061out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg062out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg063out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg064out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg065out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg066out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg067out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg068out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg069out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg070out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg071out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg072out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg073out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg074out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg075out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg076out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg077out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg078out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg079out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg080out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg081out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg082out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg083out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg084out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg085out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg086out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg087out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg088out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg089out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg090out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg091out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg092out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg093out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg094out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg095out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg096out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg097out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg098out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg099out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg100out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg101out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg102out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg103out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg104out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg105out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg106out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg107out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg108out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg109out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg110out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg111out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg112out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg113out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg114out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg115out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg116out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg117out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg118out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg119out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg120out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg121out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg122out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg123out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg124out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg125out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg126out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg127out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg128out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg129out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg130out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg131out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg132out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg133out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg134out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg135out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg136out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg137out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg138out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg139out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg140out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg141out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg142out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg143out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg144out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg145out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg146out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg147out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg148out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg149out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg150out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg151out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg152out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg153out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg154out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg155out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg156out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg157out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg158out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg159out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg160out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg161out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg162out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg163out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg164out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg165out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg166out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg167out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg168out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg169out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg170out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg171out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg172out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg173out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg174out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg175out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg176out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg177out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg178out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg179out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg180out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg181out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg182out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg183out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg184out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg185out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg186out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg187out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg188out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg189out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg190out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg191out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg192out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg193out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg194out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg195out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg196out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg197out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg198out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg199out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg200out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg201out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg202out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg203out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg204out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg205out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg206out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg207out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg208out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg209out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg210out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg211out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg212out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg213out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg214out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg215out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg216out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg217out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg218out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg219out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg220out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg221out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg222out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg223out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg224out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg225out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg226out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg227out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg228out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg229out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg230out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg231out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg232out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg233out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg234out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg235out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg236out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg237out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg238out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg239out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg240out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg241out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg242out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg243out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg244out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg245out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg246out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg247out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg248out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg249out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg250out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg251out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg252out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg253out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg254out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg255out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    reg256out   	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0)
  );
end black_white_filter_logic;

architecture IMP of black_white_filter_logic is
  
begin
  process (clk)
  begin
    if clk'event and clk = '1' then
      if (to_integer(unsigned(reg001in)) < THRESHOLD) then
		reg001out <= (others => '0');
	  else
		reg001out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg002in)) < THRESHOLD) then
		reg002out <= (others => '0');
	  else
		reg002out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg003in)) < THRESHOLD) then
		reg003out <= (others => '0');
	  else
		reg003out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg004in)) < THRESHOLD) then
		reg004out <= (others => '0');
	  else
		reg004out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg005in)) < THRESHOLD) then
		reg005out <= (others => '0');
	  else
		reg005out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg006in)) < THRESHOLD) then
		reg006out <= (others => '0');
	  else
		reg006out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg007in)) < THRESHOLD) then
		reg007out <= (others => '0');
	  else
		reg007out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg008in)) < THRESHOLD) then
		reg008out <= (others => '0');
	  else
		reg008out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg009in)) < THRESHOLD) then
		reg009out <= (others => '0');
	  else
		reg009out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg010in)) < THRESHOLD) then
		reg010out <= (others => '0');
	  else
		reg010out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg011in)) < THRESHOLD) then
		reg011out <= (others => '0');
	  else
		reg011out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg012in)) < THRESHOLD) then
		reg012out <= (others => '0');
	  else
		reg012out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg013in)) < THRESHOLD) then
		reg013out <= (others => '0');
	  else
		reg013out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg014in)) < THRESHOLD) then
		reg014out <= (others => '0');
	  else
		reg014out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg015in)) < THRESHOLD) then
		reg015out <= (others => '0');
	  else
		reg015out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg016in)) < THRESHOLD) then
		reg016out <= (others => '0');
	  else
		reg016out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg017in)) < THRESHOLD) then
		reg017out <= (others => '0');
	  else
		reg017out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg018in)) < THRESHOLD) then
		reg018out <= (others => '0');
	  else
		reg018out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg019in)) < THRESHOLD) then
		reg019out <= (others => '0');
	  else
		reg019out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg020in)) < THRESHOLD) then
		reg020out <= (others => '0');
	  else
		reg020out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg021in)) < THRESHOLD) then
		reg021out <= (others => '0');
	  else
		reg021out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg022in)) < THRESHOLD) then
		reg022out <= (others => '0');
	  else
		reg022out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg023in)) < THRESHOLD) then
		reg023out <= (others => '0');
	  else
		reg023out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg024in)) < THRESHOLD) then
		reg024out <= (others => '0');
	  else
		reg024out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg025in)) < THRESHOLD) then
		reg025out <= (others => '0');
	  else
		reg025out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg026in)) < THRESHOLD) then
		reg026out <= (others => '0');
	  else
		reg026out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg027in)) < THRESHOLD) then
		reg027out <= (others => '0');
	  else
		reg027out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg028in)) < THRESHOLD) then
		reg028out <= (others => '0');
	  else
		reg028out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg029in)) < THRESHOLD) then
		reg029out <= (others => '0');
	  else
		reg029out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg030in)) < THRESHOLD) then
		reg030out <= (others => '0');
	  else
		reg030out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg031in)) < THRESHOLD) then
		reg031out <= (others => '0');
	  else
		reg031out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg032in)) < THRESHOLD) then
		reg032out <= (others => '0');
	  else
		reg032out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg033in)) < THRESHOLD) then
		reg033out <= (others => '0');
	  else
		reg033out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg034in)) < THRESHOLD) then
		reg034out <= (others => '0');
	  else
		reg034out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg035in)) < THRESHOLD) then
		reg035out <= (others => '0');
	  else
		reg035out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg036in)) < THRESHOLD) then
		reg036out <= (others => '0');
	  else
		reg036out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg037in)) < THRESHOLD) then
		reg037out <= (others => '0');
	  else
		reg037out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg038in)) < THRESHOLD) then
		reg038out <= (others => '0');
	  else
		reg038out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg039in)) < THRESHOLD) then
		reg039out <= (others => '0');
	  else
		reg039out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg040in)) < THRESHOLD) then
		reg040out <= (others => '0');
	  else
		reg040out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg041in)) < THRESHOLD) then
		reg041out <= (others => '0');
	  else
		reg041out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg042in)) < THRESHOLD) then
		reg042out <= (others => '0');
	  else
		reg042out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg043in)) < THRESHOLD) then
		reg043out <= (others => '0');
	  else
		reg043out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg044in)) < THRESHOLD) then
		reg044out <= (others => '0');
	  else
		reg044out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg045in)) < THRESHOLD) then
		reg045out <= (others => '0');
	  else
		reg045out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg046in)) < THRESHOLD) then
		reg046out <= (others => '0');
	  else
		reg046out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg047in)) < THRESHOLD) then
		reg047out <= (others => '0');
	  else
		reg047out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg048in)) < THRESHOLD) then
		reg048out <= (others => '0');
	  else
		reg048out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg049in)) < THRESHOLD) then
		reg049out <= (others => '0');
	  else
		reg049out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg010in)) < THRESHOLD) then
		reg010out <= (others => '0');
	  else
		reg050out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg051in)) < THRESHOLD) then
		reg051out <= (others => '0');
	  else
		reg051out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg052in)) < THRESHOLD) then
		reg052out <= (others => '0');
	  else
		reg052out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg053in)) < THRESHOLD) then
		reg053out <= (others => '0');
	  else
		reg053out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg054in)) < THRESHOLD) then
		reg054out <= (others => '0');
	  else
		reg054out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg055in)) < THRESHOLD) then
		reg055out <= (others => '0');
	  else
		reg055out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg056in)) < THRESHOLD) then
		reg056out <= (others => '0');
	  else
		reg056out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg057in)) < THRESHOLD) then
		reg057out <= (others => '0');
	  else
		reg057out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg058in)) < THRESHOLD) then
		reg058out <= (others => '0');
	  else
		reg058out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg059in)) < THRESHOLD) then
		reg059out <= (others => '0');
	  else
		reg059out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg060in)) < THRESHOLD) then
		reg060out <= (others => '0');
	  else
		reg060out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg061in)) < THRESHOLD) then
		reg061out <= (others => '0');
	  else
		reg061out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg062in)) < THRESHOLD) then
		reg062out <= (others => '0');
	  else
		reg062out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg063in)) < THRESHOLD) then
		reg063out <= (others => '0');
	  else
		reg063out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg064in)) < THRESHOLD) then
		reg064out <= (others => '0');
	  else
		reg064out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg065in)) < THRESHOLD) then
		reg065out <= (others => '0');
	  else
		reg065out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg066in)) < THRESHOLD) then
		reg066out <= (others => '0');
	  else
		reg066out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg067in)) < THRESHOLD) then
		reg067out <= (others => '0');
	  else
		reg067out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg068in)) < THRESHOLD) then
		reg068out <= (others => '0');
	  else
		reg068out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg069in)) < THRESHOLD) then
		reg069out <= (others => '0');
	  else
		reg069out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg070in)) < THRESHOLD) then
		reg070out <= (others => '0');
	  else
		reg070out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg071in)) < THRESHOLD) then
		reg071out <= (others => '0');
	  else
		reg071out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg072in)) < THRESHOLD) then
		reg072out <= (others => '0');
	  else
		reg072out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg073in)) < THRESHOLD) then
		reg073out <= (others => '0');
	  else
		reg073out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg074in)) < THRESHOLD) then
		reg074out <= (others => '0');
	  else
		reg074out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg075in)) < THRESHOLD) then
		reg075out <= (others => '0');
	  else
		reg075out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg076in)) < THRESHOLD) then
		reg076out <= (others => '0');
	  else
		reg076out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg077in)) < THRESHOLD) then
		reg077out <= (others => '0');
	  else
		reg077out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg078in)) < THRESHOLD) then
		reg078out <= (others => '0');
	  else
		reg078out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg079in)) < THRESHOLD) then
		reg079out <= (others => '0');
	  else
		reg079out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg080in)) < THRESHOLD) then
		reg080out <= (others => '0');
	  else
		reg080out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg081in)) < THRESHOLD) then
		reg081out <= (others => '0');
	  else
		reg081out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg082in)) < THRESHOLD) then
		reg082out <= (others => '0');
	  else
		reg082out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg083in)) < THRESHOLD) then
		reg083out <= (others => '0');
	  else
		reg083out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg084in)) < THRESHOLD) then
		reg084out <= (others => '0');
	  else
		reg084out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg085in)) < THRESHOLD) then
		reg085out <= (others => '0');
	  else
		reg085out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg086in)) < THRESHOLD) then
		reg086out <= (others => '0');
	  else
		reg086out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg087in)) < THRESHOLD) then
		reg087out <= (others => '0');
	  else
		reg087out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg088in)) < THRESHOLD) then
		reg088out <= (others => '0');
	  else
		reg088out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg089in)) < THRESHOLD) then
		reg089out <= (others => '0');
	  else
		reg089out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg090in)) < THRESHOLD) then
		reg090out <= (others => '0');
	  else
		reg090out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg091in)) < THRESHOLD) then
		reg091out <= (others => '0');
	  else
		reg091out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg092in)) < THRESHOLD) then
		reg092out <= (others => '0');
	  else
		reg092out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg093in)) < THRESHOLD) then
		reg093out <= (others => '0');
	  else
		reg093out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg094in)) < THRESHOLD) then
		reg094out <= (others => '0');
	  else
		reg094out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg095in)) < THRESHOLD) then
		reg095out <= (others => '0');
	  else
		reg095out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg096in)) < THRESHOLD) then
		reg096out <= (others => '0');
	  else
		reg096out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg097in)) < THRESHOLD) then
		reg097out <= (others => '0');
	  else
		reg097out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg098in)) < THRESHOLD) then
		reg098out <= (others => '0');
	  else
		reg098out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg099in)) < THRESHOLD) then
		reg099out <= (others => '0');
	  else
		reg099out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg100in)) < THRESHOLD) then
		reg100out <= (others => '0');
	  else
		reg100out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg101in)) < THRESHOLD) then
		reg101out <= (others => '0');
	  else
		reg101out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg102in)) < THRESHOLD) then
		reg102out <= (others => '0');
	  else
		reg102out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg103in)) < THRESHOLD) then
		reg103out <= (others => '0');
	  else
		reg103out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg104in)) < THRESHOLD) then
		reg104out <= (others => '0');
	  else
		reg104out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg105in)) < THRESHOLD) then
		reg105out <= (others => '0');
	  else
		reg105out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg106in)) < THRESHOLD) then
		reg106out <= (others => '0');
	  else
		reg106out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg107in)) < THRESHOLD) then
		reg107out <= (others => '0');
	  else
		reg107out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg108in)) < THRESHOLD) then
		reg108out <= (others => '0');
	  else
		reg108out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg109in)) < THRESHOLD) then
		reg109out <= (others => '0');
	  else
		reg109out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg110in)) < THRESHOLD) then
		reg110out <= (others => '0');
	  else
		reg110out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg111in)) < THRESHOLD) then
		reg111out <= (others => '0');
	  else
		reg111out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg112in)) < THRESHOLD) then
		reg112out <= (others => '0');
	  else
		reg112out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg113in)) < THRESHOLD) then
		reg113out <= (others => '0');
	  else
		reg113out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg114in)) < THRESHOLD) then
		reg114out <= (others => '0');
	  else
		reg114out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg115in)) < THRESHOLD) then
		reg115out <= (others => '0');
	  else
		reg115out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg116in)) < THRESHOLD) then
		reg116out <= (others => '0');
	  else
		reg116out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg117in)) < THRESHOLD) then
		reg117out <= (others => '0');
	  else
		reg117out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg118in)) < THRESHOLD) then
		reg118out <= (others => '0');
	  else
		reg118out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg119in)) < THRESHOLD) then
		reg119out <= (others => '0');
	  else
		reg119out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg120in)) < THRESHOLD) then
		reg120out <= (others => '0');
	  else
		reg120out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg121in)) < THRESHOLD) then
		reg121out <= (others => '0');
	  else
		reg121out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg122in)) < THRESHOLD) then
		reg122out <= (others => '0');
	  else
		reg122out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg123in)) < THRESHOLD) then
		reg123out <= (others => '0');
	  else
		reg123out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg124in)) < THRESHOLD) then
		reg124out <= (others => '0');
	  else
		reg124out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg125in)) < THRESHOLD) then
		reg125out <= (others => '0');
	  else
		reg125out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg126in)) < THRESHOLD) then
		reg126out <= (others => '0');
	  else
		reg126out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg127in)) < THRESHOLD) then
		reg127out <= (others => '0');
	  else
		reg127out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg128in)) < THRESHOLD) then
		reg128out <= (others => '0');
	  else
		reg128out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg129in)) < THRESHOLD) then
		reg129out <= (others => '0');
	  else
		reg129out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg130in)) < THRESHOLD) then
		reg130out <= (others => '0');
	  else
		reg130out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg131in)) < THRESHOLD) then
		reg131out <= (others => '0');
	  else
		reg131out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg132in)) < THRESHOLD) then
		reg132out <= (others => '0');
	  else
		reg132out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg133in)) < THRESHOLD) then
		reg133out <= (others => '0');
	  else
		reg133out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg034in)) < THRESHOLD) then
		reg134out <= (others => '0');
	  else
		reg134out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg135in)) < THRESHOLD) then
		reg135out <= (others => '0');
	  else
		reg135out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg136in)) < THRESHOLD) then
		reg136out <= (others => '0');
	  else
		reg136out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg137in)) < THRESHOLD) then
		reg137out <= (others => '0');
	  else
		reg137out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg138in)) < THRESHOLD) then
		reg138out <= (others => '0');
	  else
		reg138out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg139in)) < THRESHOLD) then
		reg139out <= (others => '0');
	  else
		reg139out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg140in)) < THRESHOLD) then
		reg140out <= (others => '0');
	  else
		reg140out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg141in)) < THRESHOLD) then
		reg141out <= (others => '0');
	  else
		reg141out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg142in)) < THRESHOLD) then
		reg142out <= (others => '0');
	  else
		reg142out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg143in)) < THRESHOLD) then
		reg143out <= (others => '0');
	  else
		reg143out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg144in)) < THRESHOLD) then
		reg144out <= (others => '0');
	  else
		reg144out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg145in)) < THRESHOLD) then
		reg145out <= (others => '0');
	  else
		reg145out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg146in)) < THRESHOLD) then
		reg146out <= (others => '0');
	  else
		reg146out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg147in)) < THRESHOLD) then
		reg147out <= (others => '0');
	  else
		reg147out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg148in)) < THRESHOLD) then
		reg148out <= (others => '0');
	  else
		reg148out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg149in)) < THRESHOLD) then
		reg149out <= (others => '0');
	  else
		reg149out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg150in)) < THRESHOLD) then
		reg150out <= (others => '0');
	  else
		reg150out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg151in)) < THRESHOLD) then
		reg151out <= (others => '0');
	  else
		reg151out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg152in)) < THRESHOLD) then
		reg152out <= (others => '0');
	  else
		reg152out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg153in)) < THRESHOLD) then
		reg153out <= (others => '0');
	  else
		reg153out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg154in)) < THRESHOLD) then
		reg154out <= (others => '0');
	  else
		reg154out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg155in)) < THRESHOLD) then
		reg155out <= (others => '0');
	  else
		reg155out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg156in)) < THRESHOLD) then
		reg156out <= (others => '0');
	  else
		reg156out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg157in)) < THRESHOLD) then
		reg157out <= (others => '0');
	  else
		reg157out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg158in)) < THRESHOLD) then
		reg158out <= (others => '0');
	  else
		reg158out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg159in)) < THRESHOLD) then
		reg159out <= (others => '0');
	  else
		reg159out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg160in)) < THRESHOLD) then
		reg160out <= (others => '0');
	  else
		reg160out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg161in)) < THRESHOLD) then
		reg161out <= (others => '0');
	  else
		reg161out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg162in)) < THRESHOLD) then
		reg162out <= (others => '0');
	  else
		reg162out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg163in)) < THRESHOLD) then
		reg163out <= (others => '0');
	  else
		reg163out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg164in)) < THRESHOLD) then
		reg164out <= (others => '0');
	  else
		reg164out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg165in)) < THRESHOLD) then
		reg165out <= (others => '0');
	  else
		reg165out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg166in)) < THRESHOLD) then
		reg166out <= (others => '0');
	  else
		reg166out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg167in)) < THRESHOLD) then
		reg167out <= (others => '0');
	  else
		reg167out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg168in)) < THRESHOLD) then
		reg168out <= (others => '0');
	  else
		reg168out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg169in)) < THRESHOLD) then
		reg169out <= (others => '0');
	  else
		reg169out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg170in)) < THRESHOLD) then
		reg170out <= (others => '0');
	  else
		reg170out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg171in)) < THRESHOLD) then
		reg171out <= (others => '0');
	  else
		reg171out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg172in)) < THRESHOLD) then
		reg172out <= (others => '0');
	  else
		reg172out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg173in)) < THRESHOLD) then
		reg173out <= (others => '0');
	  else
		reg173out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg174in)) < THRESHOLD) then
		reg174out <= (others => '0');
	  else
		reg174out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg175in)) < THRESHOLD) then
		reg175out <= (others => '0');
	  else
		reg175out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg176in)) < THRESHOLD) then
		reg176out <= (others => '0');
	  else
		reg176out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg177in)) < THRESHOLD) then
		reg177out <= (others => '0');
	  else
		reg177out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg178in)) < THRESHOLD) then
		reg178out <= (others => '0');
	  else
		reg178out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg179in)) < THRESHOLD) then
		reg179out <= (others => '0');
	  else
		reg179out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg180in)) < THRESHOLD) then
		reg180out <= (others => '0');
	  else
		reg180out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg181in)) < THRESHOLD) then
		reg181out <= (others => '0');
	  else
		reg181out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg182in)) < THRESHOLD) then
		reg182out <= (others => '0');
	  else
		reg182out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg183in)) < THRESHOLD) then
		reg183out <= (others => '0');
	  else
		reg183out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg184in)) < THRESHOLD) then
		reg184out <= (others => '0');
	  else
		reg184out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg185in)) < THRESHOLD) then
		reg185out <= (others => '0');
	  else
		reg185out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg186in)) < THRESHOLD) then
		reg186out <= (others => '0');
	  else
		reg186out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg187in)) < THRESHOLD) then
		reg187out <= (others => '0');
	  else
		reg187out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg188in)) < THRESHOLD) then
		reg188out <= (others => '0');
	  else
		reg188out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg189in)) < THRESHOLD) then
		reg189out <= (others => '0');
	  else
		reg189out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg190in)) < THRESHOLD) then
		reg190out <= (others => '0');
	  else
		reg190out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg191in)) < THRESHOLD) then
		reg191out <= (others => '0');
	  else
		reg191out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg192in)) < THRESHOLD) then
		reg192out <= (others => '0');
	  else
		reg192out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg193in)) < THRESHOLD) then
		reg193out <= (others => '0');
	  else
		reg193out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg194in)) < THRESHOLD) then
		reg194out <= (others => '0');
	  else
		reg194out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg195in)) < THRESHOLD) then
		reg195out <= (others => '0');
	  else
		reg195out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg196in)) < THRESHOLD) then
		reg196out <= (others => '0');
	  else
		reg196out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg197in)) < THRESHOLD) then
		reg197out <= (others => '0');
	  else
		reg197out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg198in)) < THRESHOLD) then
		reg198out <= (others => '0');
	  else
		reg198out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg199in)) < THRESHOLD) then
		reg199out <= (others => '0');
	  else
		reg199out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg200in)) < THRESHOLD) then
		reg200out <= (others => '0');
	  else
		reg200out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg201in)) < THRESHOLD) then
		reg201out <= (others => '0');
	  else
		reg201out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg202in)) < THRESHOLD) then
		reg202out <= (others => '0');
	  else
		reg202out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg203in)) < THRESHOLD) then
		reg203out <= (others => '0');
	  else
		reg203out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg204in)) < THRESHOLD) then
		reg204out <= (others => '0');
	  else
		reg204out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg205in)) < THRESHOLD) then
		reg205out <= (others => '0');
	  else
		reg205out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg206in)) < THRESHOLD) then
		reg206out <= (others => '0');
	  else
		reg206out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg207in)) < THRESHOLD) then
		reg207out <= (others => '0');
	  else
		reg207out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg208in)) < THRESHOLD) then
		reg208out <= (others => '0');
	  else
		reg208out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg209in)) < THRESHOLD) then
		reg209out <= (others => '0');
	  else
		reg209out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg210in)) < THRESHOLD) then
		reg210out <= (others => '0');
	  else
		reg210out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg211in)) < THRESHOLD) then
		reg211out <= (others => '0');
	  else
		reg211out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg212in)) < THRESHOLD) then
		reg212out <= (others => '0');
	  else
		reg212out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg213in)) < THRESHOLD) then
		reg213out <= (others => '0');
	  else
		reg213out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg214in)) < THRESHOLD) then
		reg214out <= (others => '0');
	  else
		reg214out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg215in)) < THRESHOLD) then
		reg215out <= (others => '0');
	  else
		reg215out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg216in)) < THRESHOLD) then
		reg216out <= (others => '0');
	  else
		reg216out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg217in)) < THRESHOLD) then
		reg217out <= (others => '0');
	  else
		reg217out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg218in)) < THRESHOLD) then
		reg218out <= (others => '0');
	  else
		reg218out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg219in)) < THRESHOLD) then
		reg219out <= (others => '0');
	  else
		reg219out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg220in)) < THRESHOLD) then
		reg220out <= (others => '0');
	  else
		reg220out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg221in)) < THRESHOLD) then
		reg221out <= (others => '0');
	  else
		reg221out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg222in)) < THRESHOLD) then
		reg222out <= (others => '0');
	  else
		reg222out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg223in)) < THRESHOLD) then
		reg223out <= (others => '0');
	  else
		reg223out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg224in)) < THRESHOLD) then
		reg224out <= (others => '0');
	  else
		reg224out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg225in)) < THRESHOLD) then
		reg225out <= (others => '0');
	  else
		reg225out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg226in)) < THRESHOLD) then
		reg226out <= (others => '0');
	  else
		reg226out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg227in)) < THRESHOLD) then
		reg227out <= (others => '0');
	  else
		reg227out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg228in)) < THRESHOLD) then
		reg228out <= (others => '0');
	  else
		reg228out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg229in)) < THRESHOLD) then
		reg229out <= (others => '0');
	  else
		reg229out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg230in)) < THRESHOLD) then
		reg230out <= (others => '0');
	  else
		reg230out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg231in)) < THRESHOLD) then
		reg231out <= (others => '0');
	  else
		reg231out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg232in)) < THRESHOLD) then
		reg232out <= (others => '0');
	  else
		reg232out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg233in)) < THRESHOLD) then
		reg233out <= (others => '0');
	  else
		reg233out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg234in)) < THRESHOLD) then
		reg234out <= (others => '0');
	  else
		reg234out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg235in)) < THRESHOLD) then
		reg235out <= (others => '0');
	  else
		reg235out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg236in)) < THRESHOLD) then
		reg236out <= (others => '0');
	  else
		reg236out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg237in)) < THRESHOLD) then
		reg237out <= (others => '0');
	  else
		reg237out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg238in)) < THRESHOLD) then
		reg238out <= (others => '0');
	  else
		reg238out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg239in)) < THRESHOLD) then
		reg239out <= (others => '0');
	  else
		reg239out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg240in)) < THRESHOLD) then
		reg240out <= (others => '0');
	  else
		reg240out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg241in)) < THRESHOLD) then
		reg241out <= (others => '0');
	  else
		reg241out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg242in)) < THRESHOLD) then
		reg242out <= (others => '0');
	  else
		reg242out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg243in)) < THRESHOLD) then
		reg243out <= (others => '0');
	  else
		reg243out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg244in)) < THRESHOLD) then
		reg244out <= (others => '0');
	  else
		reg244out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg245in)) < THRESHOLD) then
		reg245out <= (others => '0');
	  else
		reg245out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg246in)) < THRESHOLD) then
		reg246out <= (others => '0');
	  else
		reg246out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg247in)) < THRESHOLD) then
		reg247out <= (others => '0');
	  else
		reg247out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg248in)) < THRESHOLD) then
		reg248out <= (others => '0');
	  else
		reg248out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg249in)) < THRESHOLD) then
		reg249out <= (others => '0');
	  else
		reg249out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg250in)) < THRESHOLD) then
		reg250out <= (others => '0');
	  else
		reg250out <= (others => '1');
	  end if;
	  if (to_integer(unsigned(reg251in)) < THRESHOLD) then
		reg251out <= (others => '0');
	  else
		reg251out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg252in)) < THRESHOLD) then
		reg252out <= (others => '0');
	  else
		reg252out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg253in)) < THRESHOLD) then
		reg253out <= (others => '0');
	  else
		reg253out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg254in)) < THRESHOLD) then
		reg254out <= (others => '0');
	  else
		reg254out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg255in)) < THRESHOLD) then
		reg255out <= (others => '0');
	  else
		reg255out <= (others => '1');
	  end if;
      if (to_integer(unsigned(reg256in)) < THRESHOLD) then
		reg256out <= (others => '0');
	  else
		reg256out <= (others => '1');
	  end if;
    end if;
  end process;
end IMP;
