-------------------------------------------------------------------------------
--
-- Top entity for testing the functionality of the top_gamma entity
--
-------------------------------------------------------------------------------
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
--
-------------------------------------------------------------------------------
--
entity top_gamma is

	-- 'clk_200MHz' are the inputs of entity.

	port (
    	clk      				: in  std_logic;
		rst						: in std_logic
	);

end top_gamma;
--
--------------------------------------------------------------------------------
--
architecture beh of top_gamma is

begin

end beh;
--
-------------------------------------------------------------------------------